`include "HardFloat/source/addRecFN.v"

module FP_Adder(
    
);


endmodule;
